`timescale 10 ns / 1 ns

`define DATA_WIDTH 32

module alu (
    input  [`DATA_WIDTH - 1:0]  A,
    input  [`DATA_WIDTH - 1:0]  B,
    input  [              2:0]  ALUop,
    output                      Overflow,
    output                      CarryOut,
    output                      Zero,
    output [`DATA_WIDTH - 1:0]  Result
);

    // Status Flags
    localparam AND = 3'b000;
    localparam  OR = 3'b001;
    localparam ADD = 3'b010;
    localparam SUB = 3'b110;
    localparam SLT = 3'b111;

    wire   [`DATA_WIDTH - 1:0]  B_trans;
    wire                        cout;
    wire   [`DATA_WIDTH - 1:0]  S;
    wire                        sign_A, sign_B, sign_S;

    // the only adder, for ADD, SUB, SLT
    adder_for_ALU alu_adder (
        .A(          A),
        .B(    B_trans),
        .cin( b_invert),
        .cout(    cout),
        .sum(        S)
    );

    // for subtraction
    assign  B_trans = {32{ALUop == SUB || ALUop == SLT}} ^ B;
    assign b_invert = ALUop == SUB || ALUop == SLT;
    // for Status Flags
    assign   sign_A = A[`DATA_WIDTH - 1];
    assign   sign_B = B[`DATA_WIDTH - 1];
    assign   sign_S = S[`DATA_WIDTH - 1];

    assign Overflow = (ALUop == ADD) & ~(sign_A ^ sign_B) & (sign_A ^ sign_S)
                    | (ALUop == SUB | ALUop == SLT) & (sign_A ^ sign_B) & (sign_A ^ sign_S);

    assign CarryOut = (ALUop == ADD) & cout
                    | (ALUop == SUB) & ((~sign_A & sign_B) | ~(sign_A ^ sign_B) & sign_S);

    assign     Zero = !Result;

    assign   Result = {32{ALUop == AND}} & (A & B)
                    | {32{ALUop == OR }} & (A | B)
                    | {32{ALUop == ADD || ALUop == SUB}} & S
                    | {32{ALUop == SLT}} & (sign_S ^ Overflow);
endmodule

module adder_for_ALU (
    input  [`DATA_WIDTH - 1:0]  A,
    input  [`DATA_WIDTH - 1:0]  B,
    input                       cin,
    output                      cout,
    output [`DATA_WIDTH - 1:0]  sum
);
    assign {cout, sum} = A + B + cin;
endmodule
